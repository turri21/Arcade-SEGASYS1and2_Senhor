localparam NOBORANKA       = 1;	// swapped address lines ($fc00 with $ff00)
localparam CHEONGCHUN      = 2;	// address and data lines swapped
localparam SHOOTING_MASTER = 3;	// light gun
localparam DAKKOCHAN       = 4; // mahjong keyboard
localparam WATER_MATCH     = 5; // special controls
